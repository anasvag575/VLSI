magic
tech scmos
timestamp 1573045415
<< rotate >>
rect 7 1 9 17
<< pwell >>
rect -6 -37 30 -14
<< nwell >>
rect -6 -1 30 22
rect 5 -5 28 -1
<< polysilicon >>
rect 1 13 3 15
rect 11 13 13 15
rect 21 13 23 15
rect 1 -24 3 3
rect 11 -24 13 3
rect 21 -24 23 3
rect 1 -30 3 -28
rect 11 -30 13 -28
rect 21 -30 23 -28
<< ndiffusion >>
rect 0 -28 1 -24
rect 3 -28 5 -24
rect 9 -28 11 -24
rect 13 -28 21 -24
rect 23 -28 24 -24
<< pdiffusion >>
rect 0 3 1 13
rect 3 3 5 13
rect 9 3 11 13
rect 13 3 15 13
rect 19 3 21 13
rect 23 3 24 13
<< metal1 >>
rect -1 17 4 21
rect 8 17 14 21
rect 18 17 24 21
rect 28 17 29 21
rect 15 13 19 17
rect -4 -17 0 3
rect 5 0 9 3
rect 24 0 28 3
rect 5 -5 28 0
rect 4 -9 9 -8
rect 14 -9 19 -8
rect 24 -9 29 -8
rect 7 -13 9 -9
rect 17 -13 19 -9
rect 27 -13 29 -9
rect 4 -14 9 -13
rect 14 -14 19 -13
rect 24 -14 29 -13
rect -4 -21 28 -17
rect 5 -24 9 -21
rect -4 -32 0 -28
rect 24 -32 28 -28
rect -5 -36 -4 -32
rect 0 -36 5 -32
rect 9 -36 15 -32
rect 19 -36 24 -32
rect 28 -36 29 -32
<< ntransistor >>
rect 1 -28 3 -24
rect 11 -28 13 -24
rect 21 -28 23 -24
<< ptransistor >>
rect 1 3 3 13
rect 11 3 13 13
rect 21 3 23 13
<< polycontact >>
rect 3 -13 7 -9
rect 13 -13 17 -9
rect 23 -13 27 -9
<< ndcontact >>
rect -4 -28 0 -24
rect 5 -28 9 -24
rect 24 -28 28 -24
<< pdcontact >>
rect -4 3 0 13
rect 5 3 9 13
rect 15 3 19 13
rect 24 3 28 13
<< psubstratepcontact >>
rect -4 -36 0 -32
rect 5 -36 9 -32
rect 15 -36 19 -32
rect 24 -36 28 -32
<< nsubstratencontact >>
rect -5 17 -1 21
rect 4 17 8 21
rect 14 17 18 21
rect 24 17 28 21
<< labels >>
rlabel metal1 29 -14 29 -8 7 C
rlabel metal1 19 -14 19 -8 1 B
rlabel metal1 9 -14 9 -8 1 A
rlabel metal1 28 -21 28 -17 7 Out
rlabel metal1 29 19 29 19 6 Vdd!
rlabel metal1 29 -34 29 -34 8 Gnd!
<< end >>
