magic
tech scmos
timestamp 1573894190
<< pwell >>
rect 121 -28 131 -24
rect -3 -40 131 -28
rect -3 -57 168 -40
rect 131 -58 168 -57
<< nwell >>
rect -3 38 168 57
rect -3 -9 131 38
rect 150 22 168 38
rect 141 -26 161 -10
<< polysilicon >>
rect 5 46 93 48
rect 5 35 7 46
rect 15 41 47 43
rect 15 35 17 41
rect 25 35 27 37
rect 35 35 37 37
rect 45 35 47 41
rect 61 40 63 46
rect 71 40 73 42
rect 81 40 83 42
rect 91 40 93 46
rect 101 40 103 42
rect 111 40 113 42
rect 121 40 123 42
rect 5 -30 7 5
rect 15 -30 17 5
rect 25 -30 27 5
rect 35 -30 37 5
rect 45 -30 47 5
rect 159 34 161 37
rect 159 5 161 24
rect 61 -30 63 0
rect 71 -30 73 0
rect 81 -30 83 0
rect 91 -30 93 0
rect 101 -30 103 0
rect 111 -30 113 0
rect 121 -30 123 0
rect 159 -2 161 1
rect 150 -14 152 -11
rect 5 -43 7 -38
rect 15 -40 17 -38
rect 25 -40 27 -38
rect 35 -43 37 -38
rect 5 -45 37 -43
rect 45 -46 47 -38
rect 150 -42 152 -24
rect 61 -44 63 -42
rect 71 -44 73 -42
rect 81 -46 83 -42
rect 91 -44 93 -42
rect 101 -44 103 -42
rect 111 -44 113 -42
rect 121 -46 123 -42
rect 45 -48 123 -46
rect 150 -49 152 -46
<< ndiffusion >>
rect 158 1 159 5
rect 161 1 162 5
rect 0 -31 5 -30
rect 4 -37 5 -31
rect 0 -38 5 -37
rect 7 -38 15 -30
rect 17 -31 25 -30
rect 17 -37 19 -31
rect 23 -37 25 -31
rect 17 -38 25 -37
rect 27 -31 35 -30
rect 27 -37 29 -31
rect 33 -37 35 -31
rect 27 -38 35 -37
rect 37 -31 45 -30
rect 37 -37 39 -31
rect 43 -37 45 -31
rect 37 -38 45 -37
rect 47 -31 52 -30
rect 47 -37 48 -31
rect 47 -38 52 -37
rect 60 -34 61 -30
rect 56 -38 61 -34
rect 60 -42 61 -38
rect 63 -42 71 -30
rect 73 -34 75 -30
rect 79 -34 81 -30
rect 73 -38 81 -34
rect 73 -42 75 -38
rect 79 -42 81 -38
rect 83 -34 85 -30
rect 89 -34 91 -30
rect 83 -38 91 -34
rect 83 -42 85 -38
rect 89 -42 91 -38
rect 93 -34 95 -30
rect 99 -34 101 -30
rect 93 -38 101 -34
rect 93 -42 95 -38
rect 99 -42 101 -38
rect 103 -34 105 -30
rect 109 -34 111 -30
rect 103 -38 111 -34
rect 103 -42 105 -38
rect 109 -42 111 -38
rect 113 -34 115 -30
rect 119 -34 121 -30
rect 113 -38 121 -34
rect 113 -42 115 -38
rect 119 -42 121 -38
rect 123 -34 124 -30
rect 123 -38 128 -34
rect 123 -42 124 -38
rect 149 -46 150 -42
rect 152 -46 153 -42
<< pdiffusion >>
rect 56 38 61 40
rect 0 34 5 35
rect 4 30 5 34
rect 0 26 5 30
rect 4 22 5 26
rect 0 18 5 22
rect 4 14 5 18
rect 0 10 5 14
rect 4 6 5 10
rect 0 5 5 6
rect 7 34 15 35
rect 7 30 9 34
rect 13 30 15 34
rect 7 26 15 30
rect 7 22 9 26
rect 13 22 15 26
rect 7 18 15 22
rect 7 14 9 18
rect 13 14 15 18
rect 7 10 15 14
rect 7 6 9 10
rect 13 6 15 10
rect 7 5 15 6
rect 17 34 25 35
rect 17 30 19 34
rect 23 30 25 34
rect 17 26 25 30
rect 17 22 19 26
rect 23 22 25 26
rect 17 18 25 22
rect 17 14 19 18
rect 23 14 25 18
rect 17 10 25 14
rect 17 6 19 10
rect 23 6 25 10
rect 17 5 25 6
rect 27 34 35 35
rect 27 30 29 34
rect 33 30 35 34
rect 27 26 35 30
rect 27 22 29 26
rect 33 22 35 26
rect 27 18 35 22
rect 27 14 29 18
rect 33 14 35 18
rect 27 10 35 14
rect 27 6 29 10
rect 33 6 35 10
rect 27 5 35 6
rect 37 5 45 35
rect 47 34 52 35
rect 47 30 48 34
rect 47 26 52 30
rect 47 22 48 26
rect 47 18 52 22
rect 47 14 48 18
rect 47 10 52 14
rect 47 6 48 10
rect 47 5 52 6
rect 60 34 61 38
rect 56 30 61 34
rect 60 26 61 30
rect 56 22 61 26
rect 60 18 61 22
rect 56 14 61 18
rect 60 10 61 14
rect 56 6 61 10
rect 60 2 61 6
rect 56 0 61 2
rect 63 38 71 40
rect 63 34 65 38
rect 69 34 71 38
rect 63 30 71 34
rect 63 26 65 30
rect 69 26 71 30
rect 63 22 71 26
rect 63 18 65 22
rect 69 18 71 22
rect 63 14 71 18
rect 63 10 65 14
rect 69 10 71 14
rect 63 6 71 10
rect 63 2 65 6
rect 69 2 71 6
rect 63 0 71 2
rect 73 38 81 40
rect 73 34 75 38
rect 79 34 81 38
rect 73 30 81 34
rect 73 26 75 30
rect 79 26 81 30
rect 73 22 81 26
rect 73 18 75 22
rect 79 18 81 22
rect 73 14 81 18
rect 73 10 75 14
rect 79 10 81 14
rect 73 6 81 10
rect 73 2 75 6
rect 79 2 81 6
rect 73 0 81 2
rect 83 0 91 40
rect 93 0 101 40
rect 103 38 111 40
rect 103 34 105 38
rect 109 34 111 38
rect 103 30 111 34
rect 103 26 105 30
rect 109 26 111 30
rect 103 22 111 26
rect 103 18 105 22
rect 109 18 111 22
rect 103 14 111 18
rect 103 10 105 14
rect 109 10 111 14
rect 103 6 111 10
rect 103 2 105 6
rect 109 2 111 6
rect 103 0 111 2
rect 113 38 121 40
rect 113 34 115 38
rect 119 34 121 38
rect 113 30 121 34
rect 113 26 115 30
rect 119 26 121 30
rect 113 22 121 26
rect 113 18 115 22
rect 119 18 121 22
rect 113 14 121 18
rect 113 10 115 14
rect 119 10 121 14
rect 113 6 121 10
rect 113 2 115 6
rect 119 2 121 6
rect 113 0 121 2
rect 123 38 128 40
rect 123 34 124 38
rect 123 30 128 34
rect 123 26 124 30
rect 123 22 128 26
rect 154 33 159 34
rect 158 25 159 33
rect 154 24 159 25
rect 161 33 166 34
rect 161 25 162 33
rect 161 24 166 25
rect 123 18 124 22
rect 123 14 128 18
rect 123 10 124 14
rect 123 6 128 10
rect 123 2 124 6
rect 123 0 128 2
rect 145 -15 150 -14
rect 149 -23 150 -15
rect 145 -24 150 -23
rect 152 -15 157 -14
rect 152 -23 153 -15
rect 152 -24 157 -23
<< metal1 >>
rect -3 51 0 55
rect 4 51 8 55
rect 12 51 16 55
rect 20 51 24 55
rect 28 51 32 55
rect 36 51 40 55
rect 44 51 48 55
rect 52 51 57 55
rect 61 51 65 55
rect 69 51 73 55
rect 77 51 81 55
rect 85 51 89 55
rect 93 51 97 55
rect 101 51 105 55
rect 109 51 113 55
rect 117 51 121 55
rect 125 51 129 55
rect 133 51 137 55
rect 141 51 145 55
rect 149 51 153 55
rect 157 51 161 55
rect 165 51 168 55
rect 0 34 4 36
rect 0 26 4 30
rect 0 18 4 22
rect 0 10 4 14
rect 0 5 4 6
rect 9 34 13 51
rect 9 26 13 30
rect 9 18 13 22
rect 9 10 13 14
rect 9 5 13 6
rect 19 34 23 36
rect 19 26 23 30
rect 19 18 23 22
rect 19 10 23 14
rect 19 5 23 6
rect 29 34 33 35
rect 29 26 33 30
rect 29 18 33 22
rect 29 10 33 14
rect 29 -8 33 6
rect 48 34 52 36
rect 48 26 52 30
rect 48 18 52 22
rect 48 10 52 14
rect 48 5 52 6
rect 56 38 60 41
rect 56 30 60 34
rect 56 22 60 26
rect 56 14 60 18
rect 56 6 60 10
rect 56 0 60 2
rect 65 38 69 51
rect 65 30 69 34
rect 65 22 69 26
rect 65 14 69 18
rect 65 6 69 10
rect 65 0 69 2
rect 75 38 79 41
rect 75 30 79 34
rect 75 22 79 26
rect 75 14 79 18
rect 75 6 79 10
rect 75 0 79 2
rect 105 38 109 40
rect 105 30 109 34
rect 105 22 109 26
rect 105 14 109 18
rect 105 6 109 10
rect 105 -3 109 2
rect 115 38 119 41
rect 115 30 119 34
rect 115 22 119 26
rect 115 14 119 18
rect 115 6 119 10
rect 115 0 119 2
rect 124 38 128 51
rect 124 30 128 34
rect 124 22 128 26
rect 124 14 128 18
rect 124 6 128 10
rect 124 0 128 2
rect 77 -7 97 -3
rect 105 -7 124 -3
rect 137 -5 141 51
rect 154 33 158 51
rect 154 24 158 25
rect 162 33 166 34
rect 162 15 166 25
rect 151 11 155 15
rect 162 11 168 15
rect 162 5 166 11
rect 154 -5 158 1
rect 47 -8 50 -7
rect 19 -11 50 -8
rect 19 -12 51 -11
rect 0 -20 1 -16
rect 10 -20 11 -16
rect 0 -31 4 -30
rect 0 -51 4 -37
rect 19 -31 23 -12
rect 31 -19 38 -15
rect 69 -19 73 -15
rect 99 -19 107 -15
rect 19 -38 23 -37
rect 29 -26 52 -22
rect 29 -31 33 -26
rect 29 -38 33 -37
rect 39 -31 43 -30
rect 39 -51 43 -37
rect 48 -31 52 -26
rect 48 -38 52 -37
rect 56 -30 60 -28
rect 85 -27 109 -23
rect 85 -30 89 -27
rect 105 -30 109 -27
rect 56 -38 60 -34
rect 75 -38 79 -34
rect 85 -38 89 -34
rect 95 -38 99 -34
rect 105 -38 109 -34
rect 115 -30 119 -7
rect 137 -9 149 -5
rect 154 -9 162 -5
rect 145 -15 149 -9
rect 145 -24 149 -23
rect 153 -15 157 -14
rect 115 -38 119 -34
rect 124 -30 128 -28
rect 153 -32 157 -23
rect 124 -38 128 -34
rect 139 -36 146 -32
rect 153 -36 168 -32
rect 153 -42 157 -36
rect 75 -51 79 -42
rect 95 -51 99 -42
rect 145 -51 149 -46
rect 162 -51 166 -46
rect -3 -55 0 -51
rect 4 -55 8 -51
rect 12 -55 16 -51
rect 20 -55 24 -51
rect 28 -55 32 -51
rect 36 -55 40 -51
rect 44 -55 48 -51
rect 52 -55 56 -51
rect 60 -55 64 -51
rect 68 -55 72 -51
rect 76 -55 80 -51
rect 84 -55 88 -51
rect 92 -55 96 -51
rect 100 -55 105 -51
rect 109 -55 113 -51
rect 117 -55 121 -51
rect 125 -55 129 -51
rect 133 -55 137 -51
rect 141 -55 145 -51
rect 149 -55 153 -51
rect 157 -55 161 -51
rect 165 -55 168 -51
<< metal2 >>
rect 60 41 75 45
rect 79 41 115 45
rect 4 36 19 40
rect 23 36 48 40
rect 134 11 147 15
rect 134 -3 138 11
rect 128 -7 138 -3
rect 54 -11 99 -7
rect 95 -15 99 -11
rect 42 -19 65 -15
rect 99 -19 139 -15
rect 60 -28 124 -24
rect 135 -32 139 -19
rect 162 -42 166 -9
<< ntransistor >>
rect 159 1 161 5
rect 5 -38 7 -30
rect 15 -38 17 -30
rect 25 -38 27 -30
rect 35 -38 37 -30
rect 45 -38 47 -30
rect 61 -42 63 -30
rect 71 -42 73 -30
rect 81 -42 83 -30
rect 91 -42 93 -30
rect 101 -42 103 -30
rect 111 -42 113 -30
rect 121 -42 123 -30
rect 150 -46 152 -42
<< ptransistor >>
rect 5 5 7 35
rect 15 5 17 35
rect 25 5 27 35
rect 35 5 37 35
rect 45 5 47 35
rect 61 0 63 40
rect 71 0 73 40
rect 81 0 83 40
rect 91 0 93 40
rect 101 0 103 40
rect 111 0 113 40
rect 121 0 123 40
rect 159 24 161 34
rect 150 -24 152 -14
<< polycontact >>
rect 1 -20 5 -16
rect 11 -20 15 -16
rect 27 -19 31 -15
rect 155 11 159 15
rect 73 -7 77 -3
rect 73 -19 77 -15
rect 97 -7 101 -3
rect 107 -19 111 -15
rect 146 -36 150 -32
<< ndcontact >>
rect 154 1 158 5
rect 162 1 166 5
rect 0 -37 4 -31
rect 19 -37 23 -31
rect 29 -37 33 -31
rect 39 -37 43 -31
rect 48 -37 52 -31
rect 56 -34 60 -30
rect 56 -42 60 -38
rect 75 -34 79 -30
rect 75 -42 79 -38
rect 85 -34 89 -30
rect 85 -42 89 -38
rect 95 -34 99 -30
rect 95 -42 99 -38
rect 105 -34 109 -30
rect 105 -42 109 -38
rect 115 -34 119 -30
rect 115 -42 119 -38
rect 124 -34 128 -30
rect 124 -42 128 -38
rect 145 -46 149 -42
rect 153 -46 157 -42
<< pdcontact >>
rect 0 30 4 34
rect 0 22 4 26
rect 0 14 4 18
rect 0 6 4 10
rect 9 30 13 34
rect 9 22 13 26
rect 9 14 13 18
rect 9 6 13 10
rect 19 30 23 34
rect 19 22 23 26
rect 19 14 23 18
rect 19 6 23 10
rect 29 30 33 34
rect 29 22 33 26
rect 29 14 33 18
rect 29 6 33 10
rect 48 30 52 34
rect 48 22 52 26
rect 48 14 52 18
rect 48 6 52 10
rect 56 34 60 38
rect 56 26 60 30
rect 56 18 60 22
rect 56 10 60 14
rect 56 2 60 6
rect 65 34 69 38
rect 65 26 69 30
rect 65 18 69 22
rect 65 10 69 14
rect 65 2 69 6
rect 75 34 79 38
rect 75 26 79 30
rect 75 18 79 22
rect 75 10 79 14
rect 75 2 79 6
rect 105 34 109 38
rect 105 26 109 30
rect 105 18 109 22
rect 105 10 109 14
rect 105 2 109 6
rect 115 34 119 38
rect 115 26 119 30
rect 115 18 119 22
rect 115 10 119 14
rect 115 2 119 6
rect 124 34 128 38
rect 124 26 128 30
rect 154 25 158 33
rect 162 25 166 33
rect 124 18 128 22
rect 124 10 128 14
rect 124 2 128 6
rect 145 -23 149 -15
rect 153 -23 157 -15
<< m2contact >>
rect 0 36 4 40
rect 56 41 60 45
rect 19 36 23 40
rect 48 36 52 40
rect 75 41 79 45
rect 115 41 119 45
rect 124 -7 128 -3
rect 147 11 151 15
rect 50 -11 54 -7
rect 38 -19 42 -15
rect 65 -19 69 -15
rect 95 -19 99 -15
rect 56 -28 60 -24
rect 162 -9 166 -5
rect 124 -28 128 -24
rect 135 -36 139 -32
rect 162 -46 166 -42
<< psubstratepcontact >>
rect 0 -55 4 -51
rect 8 -55 12 -51
rect 16 -55 20 -51
rect 24 -55 28 -51
rect 32 -55 36 -51
rect 40 -55 44 -51
rect 48 -55 52 -51
rect 56 -55 60 -51
rect 64 -55 68 -51
rect 72 -55 76 -51
rect 80 -55 84 -51
rect 88 -55 92 -51
rect 96 -55 100 -51
rect 105 -55 109 -51
rect 113 -55 117 -51
rect 121 -55 125 -51
rect 129 -55 133 -51
rect 137 -55 141 -51
rect 145 -55 149 -51
rect 153 -55 157 -51
rect 161 -55 165 -51
<< nsubstratencontact >>
rect 0 51 4 55
rect 8 51 12 55
rect 16 51 20 55
rect 24 51 28 55
rect 32 51 36 55
rect 40 51 44 55
rect 48 51 52 55
rect 57 51 61 55
rect 65 51 69 55
rect 73 51 77 55
rect 81 51 85 55
rect 89 51 93 55
rect 97 51 101 55
rect 105 51 109 55
rect 113 51 117 55
rect 121 51 125 55
rect 129 51 133 55
rect 137 51 141 55
rect 145 51 149 55
rect 153 51 157 55
rect 161 51 165 55
<< labels >>
rlabel metal1 32 -19 32 -15 1 cin
rlabel metal1 0 -20 0 -16 3 b
rlabel metal1 168 -55 168 -51 8 gnd!
rlabel metal1 168 -36 168 -32 7 cout
rlabel metal1 168 11 168 15 7 sout
rlabel metal1 168 51 168 55 6 vdd!
rlabel metal1 10 -20 10 -16 1 a
<< end >>
