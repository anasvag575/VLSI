magic
tech scmos
timestamp 1573160743
<< pwell >>
rect -6 -35 50 -20
rect -6 -36 48 -35
<< nwell >>
rect -6 -1 50 32
<< polysilicon >>
rect 11 24 43 26
rect 1 17 3 22
rect 11 17 13 24
rect 21 20 33 22
rect 21 17 23 20
rect 31 17 33 20
rect 41 17 43 24
rect 1 -23 3 2
rect 11 -23 13 2
rect 21 -23 23 2
rect 31 -23 33 2
rect 41 -23 43 2
rect 1 -29 3 -27
rect 11 -29 13 -27
rect 21 -29 23 -27
rect 31 -29 33 -27
rect 41 -29 43 -27
<< ndiffusion >>
rect 0 -27 1 -23
rect 3 -27 5 -23
rect 9 -27 11 -23
rect 13 -27 21 -23
rect 23 -27 25 -23
rect 29 -27 31 -23
rect 33 -27 35 -23
rect 39 -27 41 -23
rect 43 -27 44 -23
<< pdiffusion >>
rect 0 2 1 17
rect 3 2 5 17
rect 9 2 11 17
rect 13 2 15 17
rect 19 2 21 17
rect 23 2 25 17
rect 29 2 31 17
rect 33 2 41 17
rect 43 2 44 17
<< metal1 >>
rect -1 27 5 31
rect 9 27 14 31
rect 18 27 24 31
rect 28 27 34 31
rect 38 27 42 31
rect 46 27 49 31
rect -4 17 0 27
rect 5 20 29 24
rect 5 17 9 20
rect 25 17 29 20
rect 44 17 48 27
rect 15 -10 19 2
rect 37 -7 38 -3
rect 47 -7 48 -3
rect -4 -14 -3 -10
rect 5 -14 49 -10
rect -4 -23 0 -21
rect 5 -23 9 -14
rect 35 -23 39 -21
rect 25 -31 29 -27
rect 44 -31 48 -27
rect 0 -35 5 -31
rect 9 -35 14 -31
rect 18 -35 24 -31
rect 28 -35 32 -31
rect 36 -35 40 -31
rect 44 -35 49 -31
<< metal2 >>
rect 0 -21 35 -17
<< ntransistor >>
rect 1 -27 3 -23
rect 11 -27 13 -23
rect 21 -27 23 -23
rect 31 -27 33 -23
rect 41 -27 43 -23
<< ptransistor >>
rect 1 2 3 17
rect 11 2 13 17
rect 21 2 23 17
rect 31 2 33 17
rect 41 2 43 17
<< polycontact >>
rect -3 -14 1 -10
rect 33 -7 37 -3
rect 43 -7 47 -3
<< ndcontact >>
rect -4 -27 0 -23
rect 5 -27 9 -23
rect 25 -27 29 -23
rect 35 -27 39 -23
rect 44 -27 48 -23
<< pdcontact >>
rect -4 2 0 17
rect 5 2 9 17
rect 15 2 19 17
rect 25 2 29 17
rect 44 2 48 17
<< m2contact >>
rect -4 -21 0 -17
rect 35 -21 39 -17
<< psubstratepcontact >>
rect -4 -35 0 -31
rect 5 -35 9 -31
rect 14 -35 18 -31
rect 24 -35 28 -31
rect 32 -35 36 -31
rect 40 -35 44 -31
<< nsubstratencontact >>
rect -5 27 -1 31
rect 5 27 9 31
rect 14 27 18 31
rect 24 27 28 31
rect 34 27 38 31
rect 42 27 46 31
<< labels >>
rlabel metal1 -4 -14 -4 -10 3 B
rlabel metal1 38 -7 38 -3 1 C
rlabel metal1 48 -7 48 -3 7 A
rlabel metal1 49 27 49 31 6 Vdd!
rlabel metal1 49 -35 49 -31 8 Gnd!
rlabel metal1 49 -14 49 -10 7 Out
<< end >>
